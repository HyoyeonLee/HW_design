`timescale 1ns/1ps
module hello_world;
initial begin
$display(“\nHello World!\n”);
$finish;
end
endmodule
